@00000000
18000000
18400000
18A00000
18209100
A8210000
18600000
D8011800
9C630001
84850014
D4051814
03FFFFFC
15000000
	 
